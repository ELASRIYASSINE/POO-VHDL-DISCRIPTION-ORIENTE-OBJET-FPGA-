------PROGRAMME DIVISEUR DE FREQUENCE "EL ASRI YASSINE"------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MULTI_FREQ IS
	PORT( CLK, RST : IN STD_LOGIC;
			H1,H2: OUT STD_LOGIC
			);
END MULTI_FREQ;

ARCHITECTURE ARCH OF MULTI_FREQ is
SIGNAL CLK3Hz: INTEGER RANGE 0 TO 8333334;
SIGNAL CLK25Hz: INTEGER RANGE 0 TO 1000000;
SIGNAL W,X: STD_LOGIC;

BEGIN
-----------------PROCESS 3Hz / 333,34 msec-------------------
PROCESS(CLK,RST)
BEGIN

IF (RST = '0') THEN
	CLK3Hz <= 0;
   W <= '1';
	ELSIF (CLK'EVENT AND CLK = '1')  THEN 
   IF (CLK3Hz < 8333334) THEN CLK3Hz <= CLK3Hz+1 ;
	ELSE W <= not W;
	CLK3Hz <= 0;
	END IF;
	H1 <= W;
END IF;
END PROCESS;
-----------------PROCESS 25Hz / 40 msec-------------------
PROCESS(CLK,RST)
BEGIN
IF (RST = '0') THEN
   X <= '1';
	CLK25Hz <= 0;
	ELSIF (CLK'EVENT AND CLK = '1')  THEN 
   IF (CLK25Hz < 1000000) THEN CLK25Hz <= CLK25Hz+1 ;
	ELSE X <= not X;
	CLK25Hz <= 0;
	END IF;
	H2 <= X;

END IF;
END PROCESS;

END ARCH;




